module work7Sim;
endmodule