module m2Sim; // モジュールのシミュレーション m2
reg a; // データ入力
wire b; // 出力
clk clk1(ck); // クロック信号生成モジュールのインスタンス
m2 m2_1(a, b, ck); // モジュールのインスタンス m2
initial // シミュレーションの初期化
begin
$monitor("%b %b %b %b %b %0d",ck, a, b, m2_1.s0, m2_1.s1, $time); // モニタリング
$display("ck a b s0 s1 time") ; // ヘッダーの表示
$dumpfile("m2_re.vcd"); // 波形ファイルの指定
$dumpvars(0, m2Sim); // 波形変数の指定
a = 0; // データ入力の設定
#100 a = 1; // データ入力の設定
#100 a = 0; // データ入力の設定
#100 a = 1; // データ入力の設定
#100 a = 0; // データ入力の設定
#100 a = 1; // データ入力の設定
#100 a = 0; // データ入力の設定
#100 a = 1; // データ入力の設定
#100 a = 0; // データ入力の設定
#100 $finish;
end
endmodule
